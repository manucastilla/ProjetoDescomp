library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural :=  15;
          addrWidth: natural := 10
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin

tmp(0) := b"0000000000000000000";
tmp(1) := b"0100000000000000000";
tmp(2) := b"0100000100000000000";
tmp(3) := b"0100001000000000000";
tmp(4) := b"0100011010000000000";
tmp(5) := b"0100000110000000000";
tmp(6) := b"0100001010000000000";
tmp(7) := b"1000000000000111000";
tmp(8) := b"1000000100000100100";
tmp(9) := b"1000001000000010000";
tmp(10):= b"1000011010001000010";
tmp(11):= b"1000000110000101110";
tmp(12):= b"1000001010000011010";
tmp(13):= b"0101001110000000000";
tmp(14):= b"0011001110000000001";
tmp(15):= b"0110000000000111100";
tmp(16):= b"0101001100000010100";
tmp(17):= b"0011001100000000000";
tmp(18):= b"0110000000000000110";
tmp(19):= b"0101001100000010101";
tmp(20):= b"0011000000000001001";
tmp(21):= b"0110000000000010111";
tmp(22):= b"0000000000000000001";
tmp(23):= b"0111000000000000110";
tmp(24):= b"0100000000000000000";
tmp(25):= b"0011011010000000101";
tmp(26):= b"0110000000000011100";
tmp(27):= b"0000011010000000001";
tmp(28):= b"0111000000000000110";
tmp(29):= b"0100011010000000000";
tmp(30):= b"0011000100000001001";
tmp(31):= b"0110000000000100001";
tmp(32):= b"0000000100000000001";
tmp(33):= b"0111000000000000110";
tmp(34):= b"0100000100000000000";
tmp(35):= b"0011000110000000101";
tmp(36):= b"0110000000000100110";
tmp(37):= b"0000000110000000001";
tmp(38):= b"0111000000000000110";
tmp(39):= b"0100000110000000000";
tmp(40):= b"0011001000000001001";
tmp(41):= b"0110000000000101101";
tmp(42):= b"0011001000000000100";
tmp(43):= b"0110000000000110001";
tmp(44):= b"0000001000000000001";
tmp(45):= b"0111000000000000110";
tmp(46):= b"0100001000000000000";
tmp(47):= b"0011001010000000010";
tmp(48):= b"0000001010000000001";
tmp(49):= b"0111000000000000110";
tmp(50):= b"0011001010000000010";
tmp(51):= b"0110000000000110101";
tmp(52):= b"0000001000000000001";
tmp(53):= b"0111000000000000110";
tmp(54):= b"0100000000000000000";
tmp(55):= b"0100000100000000000";
tmp(56):= b"0100001000000000000";
tmp(57):= b"0100011010000000000";
tmp(58):= b"0100000110000000000";
tmp(59):= b"0100001010000000000";
tmp(60):= b"0111000000000000110";
tmp(61):= b"0101010010000001000";
tmp(62):= b"0010010010000000001";
tmp(63):= b"0011010010000000001";
tmp(64):= b"0011000100000001001";
tmp(65):= b"0100000100000000000";
tmp(66):= b"0000000100000000001";
tmp(67):= b"0111000000000000110";
tmp(68):= b"0101010100000001001";
tmp(69):= b"0010010100000000001";
tmp(70):= b"0011010100000000001";
tmp(71):= b"0011000110000000101";
tmp(72):= b"0100000110000000000";
tmp(73):= b"0000000110000000001";
tmp(74):= b"0111000000000000110";
tmp(75):= b"0101010110000001010";
tmp(76):= b"0010010110000000001";
tmp(77):= b"0011010110000000001";
tmp(78):= b"0011001000000000011";
tmp(79):= b"0110000000001010011";
tmp(80):= b"0011001000000001001";
tmp(81):= b"0100001000000000000";
tmp(82):= b"0000001000000000001";
tmp(83):= b"0111000000000000110";
tmp(84):= b"0011001010000000010";
tmp(85):= b"0100001000000000000";
tmp(86):= b"0111000000000001100";
tmp(87):= b"0101011000000001011";
tmp(88):= b"0010011000000000001";
tmp(89):= b"0011011000000000001";
tmp(90):= b"0011000110000000010";
tmp(91):= b"0100000110000000000";
tmp(92):= b"0000000110000000001";
tmp(93):= b"0111000000000000110";

		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;