library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural :=  15;
          addrWidth: natural := 10
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin

tmp(0):= b"0010000000000000000";
tmp(1):= b"0010000100000000000";
tmp(2):= b"0010001000000000000";
tmp(3):= b"0010011010000000000";
tmp(4):= b"0010000110000000000";
tmp(5):= b"0010001010000000000";
tmp(6):= b"0111000000000111000";
tmp(7):= b"0111000100000100100";
tmp(8):= b"0111001000000010000";
tmp(9):= b"0111011010001000010";
tmp(10):= b"0111000110000101110";
tmp(11):= b"0111001010000011010";
tmp(12):= b"0110001110000000000";
tmp(13):= b"1000001110000000001";
tmp(14):= b"0011001110000000001";
tmp(15):= b"0101000000000111101";
tmp(16):= b"0110001100001001100";
tmp(17):= b"0011001100000000000";
tmp(18):= b"0101000000000000110";
tmp(19):= b"0110001100001010110";
tmp(20):= b"0011000000000001001";
tmp(21):= b"0101000000000011000";
tmp(22):= b"0001000000000000001";
tmp(23):= b"0100000000000000110";
tmp(24):= b"0010000000000000000";
tmp(25):= b"0011011010000000101";
tmp(26):= b"0101000000000011101";
tmp(27):= b"0001011010000000001";
tmp(28):= b"0100000000000000110";
tmp(29):= b"0010011010000000000";
tmp(30):= b"0011000100000001001";
tmp(31):= b"0101000000000100010";
tmp(32):= b"0001000100000000001";
tmp(33):= b"0100000000000000110";
tmp(34):= b"0010000100000000000";
tmp(35):= b"0011000110000000101";
tmp(36):= b"0101000000000100111";
tmp(37):= b"0001000110000000001";
tmp(38):= b"0100000000000000110";
tmp(39):= b"0010000110000000000";
tmp(40):= b"0011001000000001001";
tmp(41):= b"0101000000000101110";
tmp(42):= b"0011001000000000100";
tmp(43):= b"0101000000000110010";
tmp(44):= b"0001001000000000001";
tmp(45):= b"0100000000000000110";
tmp(46):= b"0010001000000000000";
tmp(47):= b"0011001010000000010";
tmp(48):= b"0001001010000000001";
tmp(49):= b"0100000000000000110";
tmp(50):= b"0011001010000000010";
tmp(51):= b"0101000000000110110";
tmp(52):= b"0001001000000000001";
tmp(53):= b"0100000000000000110";
tmp(54):= b"0010000000000000000";
tmp(55):= b"0010000100000000000";
tmp(56):= b"0010001000000000000";
tmp(57):= b"0010011010000000000";
tmp(58):= b"0010000110000000000";
tmp(59):= b"0010001010000000000";
tmp(60):= b"0100000000000000110";
tmp(61):= b"0110010010000001000";
tmp(62):= b"0011010010000000000";
tmp(63):= b"0101000000001001010";
tmp(64):= b"0110010100000001001";
tmp(65):= b"0011010100000000000";
tmp(66):= b"0101000000001001110";
tmp(67):= b"0110010110000001010";
tmp(68):= b"0011010110000000000";
tmp(69):= b"0101000000001010010";
tmp(70):= b"0110011000000001011";
tmp(71):= b"0011011000000000000";
tmp(72):= b"0101000000001010110";
tmp(73):= b"0100000000000000110";
tmp(74):= b"0110010010000001000";
tmp(75):= b"0011010010000000001";
tmp(76):= b"0101000000000011101";
tmp(77):= b"0100000000001001010";
tmp(78):= b"0110010100000001001";
tmp(79):= b"0011010100000000001";
tmp(80):= b"0101000000000100010";
tmp(81):= b"0100000000001001110";
tmp(82):= b"0110010110000001010";
tmp(83):= b"0011010110000000001";
tmp(84):= b"0101000000000100111";
tmp(85):= b"0100000000001010010";
tmp(86):= b"0110011000000001011";
tmp(87):= b"0011011000000000001";
tmp(88):= b"0101000000000101110";
tmp(89):= b"0100000000001010110";














		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;